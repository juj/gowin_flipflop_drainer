module flipflop_drainer(
  input hdmi_clk,
  input [2:0] i_hve,
  input [23:0] i_color,
  input [12:0] x,
  input [12:0] y,
  output reg [2:0] o_hve,
  output reg [23:0] o_color
);

  reg active;
  always @(posedge hdmi_clk) begin
    o_hve <= i_hve;
    active <= (x >= 16 && y >= 16 && x < 32 && y < 32);
    o_color <= active ? {6{a449}} : i_color; // Uncomment this line to make the test case break
//    o_color <= active ? {6{a0}} : i_color; // Uncomment this line to observe the test case work
  end

  reg [3:0] a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42, a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56, a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70, a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84, a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98, a99, a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110, a111, a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122, a123, a124, a125, a126, a127, a128, a129, a130, a131, a132, a133, a134, a135, a136, a137, a138, a139, a140, a141, a142, a143, a144, a145, a146, a147, a148, a149, a150, a151, a152, a153, a154, a155, a156, a157, a158, a159, a160, a161, a162, a163, a164, a165, a166, a167, a168, a169, a170, a171, a172, a173, a174, a175, a176, a177, a178, a179, a180, a181, a182, a183, a184, a185, a186, a187, a188, a189, a190, a191, a192, a193, a194, a195, a196, a197, a198, a199, a200, a201, a202, a203, a204, a205, a206, a207, a208, a209, a210, a211, a212, a213, a214, a215, a216, a217, a218, a219, a220, a221, a222, a223, a224, a225, a226, a227, a228, a229, a230, a231, a232, a233, a234, a235, a236, a237, a238, a239, a240, a241, a242, a243, a244, a245, a246, a247, a248, a249, a250, a251, a252, a253, a254, a255, a256, a257, a258, a259, a260, a261, a262, a263, a264, a265, a266, a267, a268, a269, a270, a271, a272, a273, a274, a275, a276, a277, a278, a279, a280, a281, a282, a283, a284, a285, a286, a287, a288, a289, a290, a291, a292, a293, a294, a295, a296, a297, a298, a299, a300, a301, a302, a303, a304, a305, a306, a307, a308, a309, a310, a311, a312, a313, a314, a315, a316, a317, a318, a319, a320, a321, a322, a323, a324, a325, a326, a327, a328, a329, a330, a331, a332, a333, a334, a335, a336, a337, a338, a339, a340, a341, a342, a343, a344, a345, a346, a347, a348, a349, a350, a351, a352, a353, a354, a355, a356, a357, a358, a359, a360, a361, a362, a363, a364, a365, a366, a367, a368, a369, a370, a371, a372, a373, a374, a375, a376, a377, a378, a379, a380, a381, a382, a383, a384, a385, a386, a387, a388, a389, a390, a391, a392, a393, a394, a395, a396, a397, a398, a399, a400, a401, a402, a403, a404, a405, a406, a407, a408, a409, a410, a411, a412, a413, a414, a415, a416, a417, a418, a419, a420, a421, a422, a423, a424, a425, a426, a427, a428, a429, a430, a431, a432, a433, a434, a435, a436, a437, a438, a439, a440, a441, a442, a443, a444, a445, a446, a447, a448, a449;
  always @(posedge hdmi_clk) begin
    a0 <= a0 + 1'b1;
    a1 <= a1 + a0;
    a2 <= a2 + a1;
    a3 <= a3 + a2;
    a4 <= a4 + a3;
    a5 <= a5 + a4;
    a6 <= a6 + a5;
    a7 <= a7 + a6;
    a8 <= a8 + a7;
    a9 <= a9 + a8;
    a10 <= a10 + a9;
    a11 <= a11 + a10;
    a12 <= a12 + a11;
    a13 <= a13 + a12;
    a14 <= a14 + a13;
    a15 <= a15 + a14;
    a16 <= a16 + a15;
    a17 <= a17 + a16;
    a18 <= a18 + a17;
    a19 <= a19 + a18;
    a20 <= a20 + a19;
    a21 <= a21 + a20;
    a22 <= a22 + a21;
    a23 <= a23 + a22;
    a24 <= a24 + a23;
    a25 <= a25 + a24;
    a26 <= a26 + a25;
    a27 <= a27 + a26;
    a28 <= a28 + a27;
    a29 <= a29 + a28;
    a30 <= a30 + a29;
    a31 <= a31 + a30;
    a32 <= a32 + a31;
    a33 <= a33 + a32;
    a34 <= a34 + a33;
    a35 <= a35 + a34;
    a36 <= a36 + a35;
    a37 <= a37 + a36;
    a38 <= a38 + a37;
    a39 <= a39 + a38;
    a40 <= a40 + a39;
    a41 <= a41 + a40;
    a42 <= a42 + a41;
    a43 <= a43 + a42;
    a44 <= a44 + a43;
    a45 <= a45 + a44;
    a46 <= a46 + a45;
    a47 <= a47 + a46;
    a48 <= a48 + a47;
    a49 <= a49 + a48;
    a50 <= a50 + a49;
    a51 <= a51 + a50;
    a52 <= a52 + a51;
    a53 <= a53 + a52;
    a54 <= a54 + a53;
    a55 <= a55 + a54;
    a56 <= a56 + a55;
    a57 <= a57 + a56;
    a58 <= a58 + a57;
    a59 <= a59 + a58;
    a60 <= a60 + a59;
    a61 <= a61 + a60;
    a62 <= a62 + a61;
    a63 <= a63 + a62;
    a64 <= a64 + a63;
    a65 <= a65 + a64;
    a66 <= a66 + a65;
    a67 <= a67 + a66;
    a68 <= a68 + a67;
    a69 <= a69 + a68;
    a70 <= a70 + a69;
    a71 <= a71 + a70;
    a72 <= a72 + a71;
    a73 <= a73 + a72;
    a74 <= a74 + a73;
    a75 <= a75 + a74;
    a76 <= a76 + a75;
    a77 <= a77 + a76;
    a78 <= a78 + a77;
    a79 <= a79 + a78;
    a80 <= a80 + a79;
    a81 <= a81 + a80;
    a82 <= a82 + a81;
    a83 <= a83 + a82;
    a84 <= a84 + a83;
    a85 <= a85 + a84;
    a86 <= a86 + a85;
    a87 <= a87 + a86;
    a88 <= a88 + a87;
    a89 <= a89 + a88;
    a90 <= a90 + a89;
    a91 <= a91 + a90;
    a92 <= a92 + a91;
    a93 <= a93 + a92;
    a94 <= a94 + a93;
    a95 <= a95 + a94;
    a96 <= a96 + a95;
    a97 <= a97 + a96;
    a98 <= a98 + a97;
    a99 <= a99 + a98;
    a100 <= a100 + a99;
    a101 <= a101 + a100;
    a102 <= a102 + a101;
    a103 <= a103 + a102;
    a104 <= a104 + a103;
    a105 <= a105 + a104;
    a106 <= a106 + a105;
    a107 <= a107 + a106;
    a108 <= a108 + a107;
    a109 <= a109 + a108;
    a110 <= a110 + a109;
    a111 <= a111 + a110;
    a112 <= a112 + a111;
    a113 <= a113 + a112;
    a114 <= a114 + a113;
    a115 <= a115 + a114;
    a116 <= a116 + a115;
    a117 <= a117 + a116;
    a118 <= a118 + a117;
    a119 <= a119 + a118;
    a120 <= a120 + a119;
    a121 <= a121 + a120;
    a122 <= a122 + a121;
    a123 <= a123 + a122;
    a124 <= a124 + a123;
    a125 <= a125 + a124;
    a126 <= a126 + a125;
    a127 <= a127 + a126;
    a128 <= a128 + a127;
    a129 <= a129 + a128;
    a130 <= a130 + a129;
    a131 <= a131 + a130;
    a132 <= a132 + a131;
    a133 <= a133 + a132;
    a134 <= a134 + a133;
    a135 <= a135 + a134;
    a136 <= a136 + a135;
    a137 <= a137 + a136;
    a138 <= a138 + a137;
    a139 <= a139 + a138;
    a140 <= a140 + a139;
    a141 <= a141 + a140;
    a142 <= a142 + a141;
    a143 <= a143 + a142;
    a144 <= a144 + a143;
    a145 <= a145 + a144;
    a146 <= a146 + a145;
    a147 <= a147 + a146;
    a148 <= a148 + a147;
    a149 <= a149 + a148;
    a150 <= a150 + a149;
    a151 <= a151 + a150;
    a152 <= a152 + a151;
    a153 <= a153 + a152;
    a154 <= a154 + a153;
    a155 <= a155 + a154;
    a156 <= a156 + a155;
    a157 <= a157 + a156;
    a158 <= a158 + a157;
    a159 <= a159 + a158;
    a160 <= a160 + a159;
    a161 <= a161 + a160;
    a162 <= a162 + a161;
    a163 <= a163 + a162;
    a164 <= a164 + a163;
    a165 <= a165 + a164;
    a166 <= a166 + a165;
    a167 <= a167 + a166;
    a168 <= a168 + a167;
    a169 <= a169 + a168;
    a170 <= a170 + a169;
    a171 <= a171 + a170;
    a172 <= a172 + a171;
    a173 <= a173 + a172;
    a174 <= a174 + a173;
    a175 <= a175 + a174;
    a176 <= a176 + a175;
    a177 <= a177 + a176;
    a178 <= a178 + a177;
    a179 <= a179 + a178;
    a180 <= a180 + a179;
    a181 <= a181 + a180;
    a182 <= a182 + a181;
    a183 <= a183 + a182;
    a184 <= a184 + a183;
    a185 <= a185 + a184;
    a186 <= a186 + a185;
    a187 <= a187 + a186;
    a188 <= a188 + a187;
    a189 <= a189 + a188;
    a190 <= a190 + a189;
    a191 <= a191 + a190;
    a192 <= a192 + a191;
    a193 <= a193 + a192;
    a194 <= a194 + a193;
    a195 <= a195 + a194;
    a196 <= a196 + a195;
    a197 <= a197 + a196;
    a198 <= a198 + a197;
    a199 <= a199 + a198;
    a200 <= a200 + a199;
    a201 <= a201 + a200;
    a202 <= a202 + a201;
    a203 <= a203 + a202;
    a204 <= a204 + a203;
    a205 <= a205 + a204;
    a206 <= a206 + a205;
    a207 <= a207 + a206;
    a208 <= a208 + a207;
    a209 <= a209 + a208;
    a210 <= a210 + a209;
    a211 <= a211 + a210;
    a212 <= a212 + a211;
    a213 <= a213 + a212;
    a214 <= a214 + a213;
    a215 <= a215 + a214;
    a216 <= a216 + a215;
    a217 <= a217 + a216;
    a218 <= a218 + a217;
    a219 <= a219 + a218;
    a220 <= a220 + a219;
    a221 <= a221 + a220;
    a222 <= a222 + a221;
    a223 <= a223 + a222;
    a224 <= a224 + a223;
    a225 <= a225 + a224;
    a226 <= a226 + a225;
    a227 <= a227 + a226;
    a228 <= a228 + a227;
    a229 <= a229 + a228;
    a230 <= a230 + a229;
    a231 <= a231 + a230;
    a232 <= a232 + a231;
    a233 <= a233 + a232;
    a234 <= a234 + a233;
    a235 <= a235 + a234;
    a236 <= a236 + a235;
    a237 <= a237 + a236;
    a238 <= a238 + a237;
    a239 <= a239 + a238;
    a240 <= a240 + a239;
    a241 <= a241 + a240;
    a242 <= a242 + a241;
    a243 <= a243 + a242;
    a244 <= a244 + a243;
    a245 <= a245 + a244;
    a246 <= a246 + a245;
    a247 <= a247 + a246;
    a248 <= a248 + a247;
    a249 <= a249 + a248;
    a250 <= a250 + a249;
    a251 <= a251 + a250;
    a252 <= a252 + a251;
    a253 <= a253 + a252;
    a254 <= a254 + a253;
    a255 <= a255 + a254;
    a256 <= a256 + a255;
    a257 <= a257 + a256;
    a258 <= a258 + a257;
    a259 <= a259 + a258;
    a260 <= a260 + a259;
    a261 <= a261 + a260;
    a262 <= a262 + a261;
    a263 <= a263 + a262;
    a264 <= a264 + a263;
    a265 <= a265 + a264;
    a266 <= a266 + a265;
    a267 <= a267 + a266;
    a268 <= a268 + a267;
    a269 <= a269 + a268;
    a270 <= a270 + a269;
    a271 <= a271 + a270;
    a272 <= a272 + a271;
    a273 <= a273 + a272;
    a274 <= a274 + a273;
    a275 <= a275 + a274;
    a276 <= a276 + a275;
    a277 <= a277 + a276;
    a278 <= a278 + a277;
    a279 <= a279 + a278;
    a280 <= a280 + a279;
    a281 <= a281 + a280;
    a282 <= a282 + a281;
    a283 <= a283 + a282;
    a284 <= a284 + a283;
    a285 <= a285 + a284;
    a286 <= a286 + a285;
    a287 <= a287 + a286;
    a288 <= a288 + a287;
    a289 <= a289 + a288;
    a290 <= a290 + a289;
    a291 <= a291 + a290;
    a292 <= a292 + a291;
    a293 <= a293 + a292;
    a294 <= a294 + a293;
    a295 <= a295 + a294;
    a296 <= a296 + a295;
    a297 <= a297 + a296;
    a298 <= a298 + a297;
    a299 <= a299 + a298;
    a300 <= a300 + a299;
    a301 <= a301 + a300;
    a302 <= a302 + a301;
    a303 <= a303 + a302;
    a304 <= a304 + a303;
    a305 <= a305 + a304;
    a306 <= a306 + a305;
    a307 <= a307 + a306;
    a308 <= a308 + a307;
    a309 <= a309 + a308;
    a310 <= a310 + a309;
    a311 <= a311 + a310;
    a312 <= a312 + a311;
    a313 <= a313 + a312;
    a314 <= a314 + a313;
    a315 <= a315 + a314;
    a316 <= a316 + a315;
    a317 <= a317 + a316;
    a318 <= a318 + a317;
    a319 <= a319 + a318;
    a320 <= a320 + a319;
    a321 <= a321 + a320;
    a322 <= a322 + a321;
    a323 <= a323 + a322;
    a324 <= a324 + a323;
    a325 <= a325 + a324;
    a326 <= a326 + a325;
    a327 <= a327 + a326;
    a328 <= a328 + a327;
    a329 <= a329 + a328;
    a330 <= a330 + a329;
    a331 <= a331 + a330;
    a332 <= a332 + a331;
    a333 <= a333 + a332;
    a334 <= a334 + a333;
    a335 <= a335 + a334;
    a336 <= a336 + a335;
    a337 <= a337 + a336;
    a338 <= a338 + a337;
    a339 <= a339 + a338;
    a340 <= a340 + a339;
    a341 <= a341 + a340;
    a342 <= a342 + a341;
    a343 <= a343 + a342;
    a344 <= a344 + a343;
    a345 <= a345 + a344;
    a346 <= a346 + a345;
    a347 <= a347 + a346;
    a348 <= a348 + a347;
    a349 <= a349 + a348;
    a350 <= a350 + a349;
    a351 <= a351 + a350;
    a352 <= a352 + a351;
    a353 <= a353 + a352;
    a354 <= a354 + a353;
    a355 <= a355 + a354;
    a356 <= a356 + a355;
    a357 <= a357 + a356;
    a358 <= a358 + a357;
    a359 <= a359 + a358;
    a360 <= a360 + a359;
    a361 <= a361 + a360;
    a362 <= a362 + a361;
    a363 <= a363 + a362;
    a364 <= a364 + a363;
    a365 <= a365 + a364;
    a366 <= a366 + a365;
    a367 <= a367 + a366;
    a368 <= a368 + a367;
    a369 <= a369 + a368;
    a370 <= a370 + a369;
    a371 <= a371 + a370;
    a372 <= a372 + a371;
    a373 <= a373 + a372;
    a374 <= a374 + a373;
    a375 <= a375 + a374;
    a376 <= a376 + a375;
    a377 <= a377 + a376;
    a378 <= a378 + a377;
    a379 <= a379 + a378;
    a380 <= a380 + a379;
    a381 <= a381 + a380;
    a382 <= a382 + a381;
    a383 <= a383 + a382;
    a384 <= a384 + a383;
    a385 <= a385 + a384;
    a386 <= a386 + a385;
    a387 <= a387 + a386;
    a388 <= a388 + a387;
    a389 <= a389 + a388;
    a390 <= a390 + a389;
    a391 <= a391 + a390;
    a392 <= a392 + a391;
    a393 <= a393 + a392;
    a394 <= a394 + a393;
    a395 <= a395 + a394;
    a396 <= a396 + a395;
    a397 <= a397 + a396;
    a398 <= a398 + a397;
    a399 <= a399 + a398;
    a400 <= a400 + a399;
    a401 <= a401 + a400;
    a402 <= a402 + a401;
    a403 <= a403 + a402;
    a404 <= a404 + a403;
    a405 <= a405 + a404;
    a406 <= a406 + a405;
    a407 <= a407 + a406;
    a408 <= a408 + a407;
    a409 <= a409 + a408;
    a410 <= a410 + a409;
    a411 <= a411 + a410;
    a412 <= a412 + a411;
    a413 <= a413 + a412;
    a414 <= a414 + a413;
    a415 <= a415 + a414;
    a416 <= a416 + a415;
    a417 <= a417 + a416;
    a418 <= a418 + a417;
    a419 <= a419 + a418;
    a420 <= a420 + a419;
    a421 <= a421 + a420;
    a422 <= a422 + a421;
    a423 <= a423 + a422;
    a424 <= a424 + a423;
    a425 <= a425 + a424;
    a426 <= a426 + a425;
    a427 <= a427 + a426;
    a428 <= a428 + a427;
    a429 <= a429 + a428;
    a430 <= a430 + a429;
    a431 <= a431 + a430;
    a432 <= a432 + a431;
    a433 <= a433 + a432;
    a434 <= a434 + a433;
    a435 <= a435 + a434;
    a436 <= a436 + a435;
    a437 <= a437 + a436;
    a438 <= a438 + a437;
    a439 <= a439 + a438;
    a440 <= a440 + a439;
    a441 <= a441 + a440;
    a442 <= a442 + a441;
    a443 <= a443 + a442;
    a444 <= a444 + a443;
    a445 <= a445 + a444;
    a446 <= a446 + a445;
    a447 <= a447 + a446;
    a448 <= a448 + a447;
    a449 <= a449 + a448;
  end
endmodule
