`include "board_config.v"

module flipflop_drainer(
  input clk,
  output reg out
);
  always @(posedge clk) begin
`ifdef GW1N4
    out <= ^a450;
`endif
`ifdef GW1N9
    out <= ^a950;
`endif
`ifdef GW2A
    out <= ^a1500;
`endif

    // out <= ^a0; // Uncomment this line to observe the test case work (this optimizes away all the additions below so they won't confuse the video signal)
  end

  reg [3:0] a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42, a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56, a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70, a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84, a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98, a99, a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110, a111, a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122, a123, a124, a125, a126, a127, a128, a129, a130, a131, a132, a133, a134, a135, a136, a137, a138, a139, a140, a141, a142, a143, a144, a145, a146, a147, a148, a149, a150, a151, a152, a153, a154, a155, a156, a157, a158, a159, a160, a161, a162, a163, a164, a165, a166, a167, a168, a169, a170, a171, a172, a173, a174, a175, a176, a177, a178, a179, a180, a181, a182, a183, a184, a185, a186, a187, a188, a189, a190, a191, a192, a193, a194, a195, a196, a197, a198, a199, a200, a201, a202, a203, a204, a205, a206, a207, a208, a209, a210, a211, a212, a213, a214, a215, a216, a217, a218, a219, a220, a221, a222, a223, a224, a225, a226, a227, a228, a229, a230, a231, a232, a233, a234, a235, a236, a237, a238, a239, a240, a241, a242, a243, a244, a245, a246, a247, a248, a249, a250, a251, a252, a253, a254, a255, a256, a257, a258, a259, a260, a261, a262, a263, a264, a265, a266, a267, a268, a269, a270, a271, a272, a273, a274, a275, a276, a277, a278, a279, a280, a281, a282, a283, a284, a285, a286, a287, a288, a289, a290, a291, a292, a293, a294, a295, a296, a297, a298, a299, a300, a301, a302, a303, a304, a305, a306, a307, a308, a309, a310, a311, a312, a313, a314, a315, a316, a317, a318, a319, a320, a321, a322, a323, a324, a325, a326, a327, a328, a329, a330, a331, a332, a333, a334, a335, a336, a337, a338, a339, a340, a341, a342, a343, a344, a345, a346, a347, a348, a349, a350, a351, a352, a353, a354, a355, a356, a357, a358, a359, a360, a361, a362, a363, a364, a365, a366, a367, a368, a369, a370, a371, a372, a373, a374, a375, a376, a377, a378, a379, a380, a381, a382, a383, a384, a385, a386, a387, a388, a389, a390, a391, a392, a393, a394, a395, a396, a397, a398, a399, a400, a401, a402, a403, a404, a405, a406, a407, a408, a409, a410, a411, a412, a413, a414, a415, a416, a417, a418, a419, a420, a421, a422, a423, a424, a425, a426, a427, a428, a429, a430, a431, a432, a433, a434, a435, a436, a437, a438, a439, a440, a441, a442, a443, a444, a445, a446, a447, a448, a449, a450, a451, a452, a453, a454, a455, a456, a457, a458, a459, a460, a461, a462, a463, a464, a465, a466, a467, a468, a469, a470, a471, a472, a473, a474, a475, a476, a477, a478, a479, a480, a481, a482, a483, a484, a485, a486, a487, a488, a489, a490, a491, a492, a493, a494, a495, a496, a497, a498, a499, a500, a501, a502, a503, a504, a505, a506, a507, a508, a509, a510, a511, a512, a513, a514, a515, a516, a517, a518, a519, a520, a521, a522, a523, a524, a525, a526, a527, a528, a529, a530, a531, a532, a533, a534, a535, a536, a537, a538, a539, a540, a541, a542, a543, a544, a545, a546, a547, a548, a549, a550, a551, a552, a553, a554, a555, a556, a557, a558, a559, a560, a561, a562, a563, a564, a565, a566, a567, a568, a569, a570, a571, a572, a573, a574, a575, a576, a577, a578, a579, a580, a581, a582, a583, a584, a585, a586, a587, a588, a589, a590, a591, a592, a593, a594, a595, a596, a597, a598, a599, a600, a601, a602, a603, a604, a605, a606, a607, a608, a609, a610, a611, a612, a613, a614, a615, a616, a617, a618, a619, a620, a621, a622, a623, a624, a625, a626, a627, a628, a629, a630, a631, a632, a633, a634, a635, a636, a637, a638, a639, a640, a641, a642, a643, a644, a645, a646, a647, a648, a649, a650, a651, a652, a653, a654, a655, a656, a657, a658, a659, a660, a661, a662, a663, a664, a665, a666, a667, a668, a669, a670, a671, a672, a673, a674, a675, a676, a677, a678, a679, a680, a681, a682, a683, a684, a685, a686, a687, a688, a689, a690, a691, a692, a693, a694, a695, a696, a697, a698, a699, a700, a701, a702, a703, a704, a705, a706, a707, a708, a709, a710, a711, a712, a713, a714, a715, a716, a717, a718, a719, a720, a721, a722, a723, a724, a725, a726, a727, a728, a729, a730, a731, a732, a733, a734, a735, a736, a737, a738, a739, a740, a741, a742, a743, a744, a745, a746, a747, a748, a749, a750, a751, a752, a753, a754, a755, a756, a757, a758, a759, a760, a761, a762, a763, a764, a765, a766, a767, a768, a769, a770, a771, a772, a773, a774, a775, a776, a777, a778, a779, a780, a781, a782, a783, a784, a785, a786, a787, a788, a789, a790, a791, a792, a793, a794, a795, a796, a797, a798, a799, a800, a801, a802, a803, a804, a805, a806, a807, a808, a809, a810, a811, a812, a813, a814, a815, a816, a817, a818, a819, a820, a821, a822, a823, a824, a825, a826, a827, a828, a829, a830, a831, a832, a833, a834, a835, a836, a837, a838, a839, a840, a841, a842, a843, a844, a845, a846, a847, a848, a849, a850, a851, a852, a853, a854, a855, a856, a857, a858, a859, a860, a861, a862, a863, a864, a865, a866, a867, a868, a869, a870, a871, a872, a873, a874, a875, a876, a877, a878, a879, a880, a881, a882, a883, a884, a885, a886, a887, a888, a889, a890, a891, a892, a893, a894, a895, a896, a897, a898, a899, a900, a901, a902, a903, a904, a905, a906, a907, a908, a909, a910, a911, a912, a913, a914, a915, a916, a917, a918, a919, a920, a921, a922, a923, a924, a925, a926, a927, a928, a929, a930, a931, a932, a933, a934, a935, a936, a937, a938, a939, a940, a941, a942, a943, a944, a945, a946, a947, a948, a949, a950, a951, a952, a953, a954, a955, a956, a957, a958, a959, a960, a961, a962, a963, a964, a965, a966, a967, a968, a969, a970, a971, a972, a973, a974, a975, a976, a977, a978, a979, a980, a981, a982, a983, a984, a985, a986, a987, a988, a989, a990, a991, a992, a993, a994, a995, a996, a997, a998, a999, a1000, a1001, a1002, a1003, a1004, a1005, a1006, a1007, a1008, a1009, a1010, a1011, a1012, a1013, a1014, a1015, a1016, a1017, a1018, a1019, a1020, a1021, a1022, a1023, a1024, a1025, a1026, a1027, a1028, a1029, a1030, a1031, a1032, a1033, a1034, a1035, a1036, a1037, a1038, a1039, a1040, a1041, a1042, a1043, a1044, a1045, a1046, a1047, a1048, a1049, a1050, a1051, a1052, a1053, a1054, a1055, a1056, a1057, a1058, a1059, a1060, a1061, a1062, a1063, a1064, a1065, a1066, a1067, a1068, a1069, a1070, a1071, a1072, a1073, a1074, a1075, a1076, a1077, a1078, a1079, a1080, a1081, a1082, a1083, a1084, a1085, a1086, a1087, a1088, a1089, a1090, a1091, a1092, a1093, a1094, a1095, a1096, a1097, a1098, a1099, a1100, a1101, a1102, a1103, a1104, a1105, a1106, a1107, a1108, a1109, a1110, a1111, a1112, a1113, a1114, a1115, a1116, a1117, a1118, a1119, a1120, a1121, a1122, a1123, a1124, a1125, a1126, a1127, a1128, a1129, a1130, a1131, a1132, a1133, a1134, a1135, a1136, a1137, a1138, a1139, a1140, a1141, a1142, a1143, a1144, a1145, a1146, a1147, a1148, a1149, a1150, a1151, a1152, a1153, a1154, a1155, a1156, a1157, a1158, a1159, a1160, a1161, a1162, a1163, a1164, a1165, a1166, a1167, a1168, a1169, a1170, a1171, a1172, a1173, a1174, a1175, a1176, a1177, a1178, a1179, a1180, a1181, a1182, a1183, a1184, a1185, a1186, a1187, a1188, a1189, a1190, a1191, a1192, a1193, a1194, a1195, a1196, a1197, a1198, a1199, a1200, a1201, a1202, a1203, a1204, a1205, a1206, a1207, a1208, a1209, a1210, a1211, a1212, a1213, a1214, a1215, a1216, a1217, a1218, a1219, a1220, a1221, a1222, a1223, a1224, a1225, a1226, a1227, a1228, a1229, a1230, a1231, a1232, a1233, a1234, a1235, a1236, a1237, a1238, a1239, a1240, a1241, a1242, a1243, a1244, a1245, a1246, a1247, a1248, a1249, a1250, a1251, a1252, a1253, a1254, a1255, a1256, a1257, a1258, a1259, a1260, a1261, a1262, a1263, a1264, a1265, a1266, a1267, a1268, a1269, a1270, a1271, a1272, a1273, a1274, a1275, a1276, a1277, a1278, a1279, a1280, a1281, a1282, a1283, a1284, a1285, a1286, a1287, a1288, a1289, a1290, a1291, a1292, a1293, a1294, a1295, a1296, a1297, a1298, a1299, a1300, a1301, a1302, a1303, a1304, a1305, a1306, a1307, a1308, a1309, a1310, a1311, a1312, a1313, a1314, a1315, a1316, a1317, a1318, a1319, a1320, a1321, a1322, a1323, a1324, a1325, a1326, a1327, a1328, a1329, a1330, a1331, a1332, a1333, a1334, a1335, a1336, a1337, a1338, a1339, a1340, a1341, a1342, a1343, a1344, a1345, a1346, a1347, a1348, a1349, a1350, a1351, a1352, a1353, a1354, a1355, a1356, a1357, a1358, a1359, a1360, a1361, a1362, a1363, a1364, a1365, a1366, a1367, a1368, a1369, a1370, a1371, a1372, a1373, a1374, a1375, a1376, a1377, a1378, a1379, a1380, a1381, a1382, a1383, a1384, a1385, a1386, a1387, a1388, a1389, a1390, a1391, a1392, a1393, a1394, a1395, a1396, a1397, a1398, a1399, a1400, a1401, a1402, a1403, a1404, a1405, a1406, a1407, a1408, a1409, a1410, a1411, a1412, a1413, a1414, a1415, a1416, a1417, a1418, a1419, a1420, a1421, a1422, a1423, a1424, a1425, a1426, a1427, a1428, a1429, a1430, a1431, a1432, a1433, a1434, a1435, a1436, a1437, a1438, a1439, a1440, a1441, a1442, a1443, a1444, a1445, a1446, a1447, a1448, a1449, a1450, a1451, a1452, a1453, a1454, a1455, a1456, a1457, a1458, a1459, a1460, a1461, a1462, a1463, a1464, a1465, a1466, a1467, a1468, a1469, a1470, a1471, a1472, a1473, a1474, a1475, a1476, a1477, a1478, a1479, a1480, a1481, a1482, a1483, a1484, a1485, a1486, a1487, a1488, a1489, a1490, a1491, a1492, a1493, a1494, a1495, a1496, a1497, a1498, a1499, a1500;
  always @(posedge clk) begin
    a0 <= a0 + 1'b1;
    a1 <= a1 + a0;
    a2 <= a2 + a1;
    a3 <= a3 + a2;
    a4 <= a4 + a3;
    a5 <= a5 + a4;
    a6 <= a6 + a5;
    a7 <= a7 + a6;
    a8 <= a8 + a7;
    a9 <= a9 + a8;
    a10 <= a10 + a9;
    a11 <= a11 + a10;
    a12 <= a12 + a11;
    a13 <= a13 + a12;
    a14 <= a14 + a13;
    a15 <= a15 + a14;
    a16 <= a16 + a15;
    a17 <= a17 + a16;
    a18 <= a18 + a17;
    a19 <= a19 + a18;
    a20 <= a20 + a19;
    a21 <= a21 + a20;
    a22 <= a22 + a21;
    a23 <= a23 + a22;
    a24 <= a24 + a23;
    a25 <= a25 + a24;
    a26 <= a26 + a25;
    a27 <= a27 + a26;
    a28 <= a28 + a27;
    a29 <= a29 + a28;
    a30 <= a30 + a29;
    a31 <= a31 + a30;
    a32 <= a32 + a31;
    a33 <= a33 + a32;
    a34 <= a34 + a33;
    a35 <= a35 + a34;
    a36 <= a36 + a35;
    a37 <= a37 + a36;
    a38 <= a38 + a37;
    a39 <= a39 + a38;
    a40 <= a40 + a39;
    a41 <= a41 + a40;
    a42 <= a42 + a41;
    a43 <= a43 + a42;
    a44 <= a44 + a43;
    a45 <= a45 + a44;
    a46 <= a46 + a45;
    a47 <= a47 + a46;
    a48 <= a48 + a47;
    a49 <= a49 + a48;
    a50 <= a50 + a49;
    a51 <= a51 + a50;
    a52 <= a52 + a51;
    a53 <= a53 + a52;
    a54 <= a54 + a53;
    a55 <= a55 + a54;
    a56 <= a56 + a55;
    a57 <= a57 + a56;
    a58 <= a58 + a57;
    a59 <= a59 + a58;
    a60 <= a60 + a59;
    a61 <= a61 + a60;
    a62 <= a62 + a61;
    a63 <= a63 + a62;
    a64 <= a64 + a63;
    a65 <= a65 + a64;
    a66 <= a66 + a65;
    a67 <= a67 + a66;
    a68 <= a68 + a67;
    a69 <= a69 + a68;
    a70 <= a70 + a69;
    a71 <= a71 + a70;
    a72 <= a72 + a71;
    a73 <= a73 + a72;
    a74 <= a74 + a73;
    a75 <= a75 + a74;
    a76 <= a76 + a75;
    a77 <= a77 + a76;
    a78 <= a78 + a77;
    a79 <= a79 + a78;
    a80 <= a80 + a79;
    a81 <= a81 + a80;
    a82 <= a82 + a81;
    a83 <= a83 + a82;
    a84 <= a84 + a83;
    a85 <= a85 + a84;
    a86 <= a86 + a85;
    a87 <= a87 + a86;
    a88 <= a88 + a87;
    a89 <= a89 + a88;
    a90 <= a90 + a89;
    a91 <= a91 + a90;
    a92 <= a92 + a91;
    a93 <= a93 + a92;
    a94 <= a94 + a93;
    a95 <= a95 + a94;
    a96 <= a96 + a95;
    a97 <= a97 + a96;
    a98 <= a98 + a97;
    a99 <= a99 + a98;
    a100 <= a100 + a99;
    a101 <= a101 + a100;
    a102 <= a102 + a101;
    a103 <= a103 + a102;
    a104 <= a104 + a103;
    a105 <= a105 + a104;
    a106 <= a106 + a105;
    a107 <= a107 + a106;
    a108 <= a108 + a107;
    a109 <= a109 + a108;
    a110 <= a110 + a109;
    a111 <= a111 + a110;
    a112 <= a112 + a111;
    a113 <= a113 + a112;
    a114 <= a114 + a113;
    a115 <= a115 + a114;
    a116 <= a116 + a115;
    a117 <= a117 + a116;
    a118 <= a118 + a117;
    a119 <= a119 + a118;
    a120 <= a120 + a119;
    a121 <= a121 + a120;
    a122 <= a122 + a121;
    a123 <= a123 + a122;
    a124 <= a124 + a123;
    a125 <= a125 + a124;
    a126 <= a126 + a125;
    a127 <= a127 + a126;
    a128 <= a128 + a127;
    a129 <= a129 + a128;
    a130 <= a130 + a129;
    a131 <= a131 + a130;
    a132 <= a132 + a131;
    a133 <= a133 + a132;
    a134 <= a134 + a133;
    a135 <= a135 + a134;
    a136 <= a136 + a135;
    a137 <= a137 + a136;
    a138 <= a138 + a137;
    a139 <= a139 + a138;
    a140 <= a140 + a139;
    a141 <= a141 + a140;
    a142 <= a142 + a141;
    a143 <= a143 + a142;
    a144 <= a144 + a143;
    a145 <= a145 + a144;
    a146 <= a146 + a145;
    a147 <= a147 + a146;
    a148 <= a148 + a147;
    a149 <= a149 + a148;
    a150 <= a150 + a149;
    a151 <= a151 + a150;
    a152 <= a152 + a151;
    a153 <= a153 + a152;
    a154 <= a154 + a153;
    a155 <= a155 + a154;
    a156 <= a156 + a155;
    a157 <= a157 + a156;
    a158 <= a158 + a157;
    a159 <= a159 + a158;
    a160 <= a160 + a159;
    a161 <= a161 + a160;
    a162 <= a162 + a161;
    a163 <= a163 + a162;
    a164 <= a164 + a163;
    a165 <= a165 + a164;
    a166 <= a166 + a165;
    a167 <= a167 + a166;
    a168 <= a168 + a167;
    a169 <= a169 + a168;
    a170 <= a170 + a169;
    a171 <= a171 + a170;
    a172 <= a172 + a171;
    a173 <= a173 + a172;
    a174 <= a174 + a173;
    a175 <= a175 + a174;
    a176 <= a176 + a175;
    a177 <= a177 + a176;
    a178 <= a178 + a177;
    a179 <= a179 + a178;
    a180 <= a180 + a179;
    a181 <= a181 + a180;
    a182 <= a182 + a181;
    a183 <= a183 + a182;
    a184 <= a184 + a183;
    a185 <= a185 + a184;
    a186 <= a186 + a185;
    a187 <= a187 + a186;
    a188 <= a188 + a187;
    a189 <= a189 + a188;
    a190 <= a190 + a189;
    a191 <= a191 + a190;
    a192 <= a192 + a191;
    a193 <= a193 + a192;
    a194 <= a194 + a193;
    a195 <= a195 + a194;
    a196 <= a196 + a195;
    a197 <= a197 + a196;
    a198 <= a198 + a197;
    a199 <= a199 + a198;
    a200 <= a200 + a199;
    a201 <= a201 + a200;
    a202 <= a202 + a201;
    a203 <= a203 + a202;
    a204 <= a204 + a203;
    a205 <= a205 + a204;
    a206 <= a206 + a205;
    a207 <= a207 + a206;
    a208 <= a208 + a207;
    a209 <= a209 + a208;
    a210 <= a210 + a209;
    a211 <= a211 + a210;
    a212 <= a212 + a211;
    a213 <= a213 + a212;
    a214 <= a214 + a213;
    a215 <= a215 + a214;
    a216 <= a216 + a215;
    a217 <= a217 + a216;
    a218 <= a218 + a217;
    a219 <= a219 + a218;
    a220 <= a220 + a219;
    a221 <= a221 + a220;
    a222 <= a222 + a221;
    a223 <= a223 + a222;
    a224 <= a224 + a223;
    a225 <= a225 + a224;
    a226 <= a226 + a225;
    a227 <= a227 + a226;
    a228 <= a228 + a227;
    a229 <= a229 + a228;
    a230 <= a230 + a229;
    a231 <= a231 + a230;
    a232 <= a232 + a231;
    a233 <= a233 + a232;
    a234 <= a234 + a233;
    a235 <= a235 + a234;
    a236 <= a236 + a235;
    a237 <= a237 + a236;
    a238 <= a238 + a237;
    a239 <= a239 + a238;
    a240 <= a240 + a239;
    a241 <= a241 + a240;
    a242 <= a242 + a241;
    a243 <= a243 + a242;
    a244 <= a244 + a243;
    a245 <= a245 + a244;
    a246 <= a246 + a245;
    a247 <= a247 + a246;
    a248 <= a248 + a247;
    a249 <= a249 + a248;
    a250 <= a250 + a249;
    a251 <= a251 + a250;
    a252 <= a252 + a251;
    a253 <= a253 + a252;
    a254 <= a254 + a253;
    a255 <= a255 + a254;
    a256 <= a256 + a255;
    a257 <= a257 + a256;
    a258 <= a258 + a257;
    a259 <= a259 + a258;
    a260 <= a260 + a259;
    a261 <= a261 + a260;
    a262 <= a262 + a261;
    a263 <= a263 + a262;
    a264 <= a264 + a263;
    a265 <= a265 + a264;
    a266 <= a266 + a265;
    a267 <= a267 + a266;
    a268 <= a268 + a267;
    a269 <= a269 + a268;
    a270 <= a270 + a269;
    a271 <= a271 + a270;
    a272 <= a272 + a271;
    a273 <= a273 + a272;
    a274 <= a274 + a273;
    a275 <= a275 + a274;
    a276 <= a276 + a275;
    a277 <= a277 + a276;
    a278 <= a278 + a277;
    a279 <= a279 + a278;
    a280 <= a280 + a279;
    a281 <= a281 + a280;
    a282 <= a282 + a281;
    a283 <= a283 + a282;
    a284 <= a284 + a283;
    a285 <= a285 + a284;
    a286 <= a286 + a285;
    a287 <= a287 + a286;
    a288 <= a288 + a287;
    a289 <= a289 + a288;
    a290 <= a290 + a289;
    a291 <= a291 + a290;
    a292 <= a292 + a291;
    a293 <= a293 + a292;
    a294 <= a294 + a293;
    a295 <= a295 + a294;
    a296 <= a296 + a295;
    a297 <= a297 + a296;
    a298 <= a298 + a297;
    a299 <= a299 + a298;
    a300 <= a300 + a299;
    a301 <= a301 + a300;
    a302 <= a302 + a301;
    a303 <= a303 + a302;
    a304 <= a304 + a303;
    a305 <= a305 + a304;
    a306 <= a306 + a305;
    a307 <= a307 + a306;
    a308 <= a308 + a307;
    a309 <= a309 + a308;
    a310 <= a310 + a309;
    a311 <= a311 + a310;
    a312 <= a312 + a311;
    a313 <= a313 + a312;
    a314 <= a314 + a313;
    a315 <= a315 + a314;
    a316 <= a316 + a315;
    a317 <= a317 + a316;
    a318 <= a318 + a317;
    a319 <= a319 + a318;
    a320 <= a320 + a319;
    a321 <= a321 + a320;
    a322 <= a322 + a321;
    a323 <= a323 + a322;
    a324 <= a324 + a323;
    a325 <= a325 + a324;
    a326 <= a326 + a325;
    a327 <= a327 + a326;
    a328 <= a328 + a327;
    a329 <= a329 + a328;
    a330 <= a330 + a329;
    a331 <= a331 + a330;
    a332 <= a332 + a331;
    a333 <= a333 + a332;
    a334 <= a334 + a333;
    a335 <= a335 + a334;
    a336 <= a336 + a335;
    a337 <= a337 + a336;
    a338 <= a338 + a337;
    a339 <= a339 + a338;
    a340 <= a340 + a339;
    a341 <= a341 + a340;
    a342 <= a342 + a341;
    a343 <= a343 + a342;
    a344 <= a344 + a343;
    a345 <= a345 + a344;
    a346 <= a346 + a345;
    a347 <= a347 + a346;
    a348 <= a348 + a347;
    a349 <= a349 + a348;
    a350 <= a350 + a349;
    a351 <= a351 + a350;
    a352 <= a352 + a351;
    a353 <= a353 + a352;
    a354 <= a354 + a353;
    a355 <= a355 + a354;
    a356 <= a356 + a355;
    a357 <= a357 + a356;
    a358 <= a358 + a357;
    a359 <= a359 + a358;
    a360 <= a360 + a359;
    a361 <= a361 + a360;
    a362 <= a362 + a361;
    a363 <= a363 + a362;
    a364 <= a364 + a363;
    a365 <= a365 + a364;
    a366 <= a366 + a365;
    a367 <= a367 + a366;
    a368 <= a368 + a367;
    a369 <= a369 + a368;
    a370 <= a370 + a369;
    a371 <= a371 + a370;
    a372 <= a372 + a371;
    a373 <= a373 + a372;
    a374 <= a374 + a373;
    a375 <= a375 + a374;
    a376 <= a376 + a375;
    a377 <= a377 + a376;
    a378 <= a378 + a377;
    a379 <= a379 + a378;
    a380 <= a380 + a379;
    a381 <= a381 + a380;
    a382 <= a382 + a381;
    a383 <= a383 + a382;
    a384 <= a384 + a383;
    a385 <= a385 + a384;
    a386 <= a386 + a385;
    a387 <= a387 + a386;
    a388 <= a388 + a387;
    a389 <= a389 + a388;
    a390 <= a390 + a389;
    a391 <= a391 + a390;
    a392 <= a392 + a391;
    a393 <= a393 + a392;
    a394 <= a394 + a393;
    a395 <= a395 + a394;
    a396 <= a396 + a395;
    a397 <= a397 + a396;
    a398 <= a398 + a397;
    a399 <= a399 + a398;
    a400 <= a400 + a399;
    a401 <= a401 + a400;
    a402 <= a402 + a401;
    a403 <= a403 + a402;
    a404 <= a404 + a403;
    a405 <= a405 + a404;
    a406 <= a406 + a405;
    a407 <= a407 + a406;
    a408 <= a408 + a407;
    a409 <= a409 + a408;
    a410 <= a410 + a409;
    a411 <= a411 + a410;
    a412 <= a412 + a411;
    a413 <= a413 + a412;
    a414 <= a414 + a413;
    a415 <= a415 + a414;
    a416 <= a416 + a415;
    a417 <= a417 + a416;
    a418 <= a418 + a417;
    a419 <= a419 + a418;
    a420 <= a420 + a419;
    a421 <= a421 + a420;
    a422 <= a422 + a421;
    a423 <= a423 + a422;
    a424 <= a424 + a423;
    a425 <= a425 + a424;
    a426 <= a426 + a425;
    a427 <= a427 + a426;
    a428 <= a428 + a427;
    a429 <= a429 + a428;
    a430 <= a430 + a429;
    a431 <= a431 + a430;
    a432 <= a432 + a431;
    a433 <= a433 + a432;
    a434 <= a434 + a433;
    a435 <= a435 + a434;
    a436 <= a436 + a435;
    a437 <= a437 + a436;
    a438 <= a438 + a437;
    a439 <= a439 + a438;
    a440 <= a440 + a439;
    a441 <= a441 + a440;
    a442 <= a442 + a441;
    a443 <= a443 + a442;
    a444 <= a444 + a443;
    a445 <= a445 + a444;
    a446 <= a446 + a445;
    a447 <= a447 + a446;
    a448 <= a448 + a447;
    a449 <= a449 + a448;
    a450 <= a450 + a449;
    a451 <= a451 + a450;
    a452 <= a452 + a451;
    a453 <= a453 + a452;
    a454 <= a454 + a453;
    a455 <= a455 + a454;
    a456 <= a456 + a455;
    a457 <= a457 + a456;
    a458 <= a458 + a457;
    a459 <= a459 + a458;
    a460 <= a460 + a459;
    a461 <= a461 + a460;
    a462 <= a462 + a461;
    a463 <= a463 + a462;
    a464 <= a464 + a463;
    a465 <= a465 + a464;
    a466 <= a466 + a465;
    a467 <= a467 + a466;
    a468 <= a468 + a467;
    a469 <= a469 + a468;
    a470 <= a470 + a469;
    a471 <= a471 + a470;
    a472 <= a472 + a471;
    a473 <= a473 + a472;
    a474 <= a474 + a473;
    a475 <= a475 + a474;
    a476 <= a476 + a475;
    a477 <= a477 + a476;
    a478 <= a478 + a477;
    a479 <= a479 + a478;
    a480 <= a480 + a479;
    a481 <= a481 + a480;
    a482 <= a482 + a481;
    a483 <= a483 + a482;
    a484 <= a484 + a483;
    a485 <= a485 + a484;
    a486 <= a486 + a485;
    a487 <= a487 + a486;
    a488 <= a488 + a487;
    a489 <= a489 + a488;
    a490 <= a490 + a489;
    a491 <= a491 + a490;
    a492 <= a492 + a491;
    a493 <= a493 + a492;
    a494 <= a494 + a493;
    a495 <= a495 + a494;
    a496 <= a496 + a495;
    a497 <= a497 + a496;
    a498 <= a498 + a497;
    a499 <= a499 + a498;
    a500 <= a500 + a499;
    a501 <= a501 + a500;
    a502 <= a502 + a501;
    a503 <= a503 + a502;
    a504 <= a504 + a503;
    a505 <= a505 + a504;
    a506 <= a506 + a505;
    a507 <= a507 + a506;
    a508 <= a508 + a507;
    a509 <= a509 + a508;
    a510 <= a510 + a509;
    a511 <= a511 + a510;
    a512 <= a512 + a511;
    a513 <= a513 + a512;
    a514 <= a514 + a513;
    a515 <= a515 + a514;
    a516 <= a516 + a515;
    a517 <= a517 + a516;
    a518 <= a518 + a517;
    a519 <= a519 + a518;
    a520 <= a520 + a519;
    a521 <= a521 + a520;
    a522 <= a522 + a521;
    a523 <= a523 + a522;
    a524 <= a524 + a523;
    a525 <= a525 + a524;
    a526 <= a526 + a525;
    a527 <= a527 + a526;
    a528 <= a528 + a527;
    a529 <= a529 + a528;
    a530 <= a530 + a529;
    a531 <= a531 + a530;
    a532 <= a532 + a531;
    a533 <= a533 + a532;
    a534 <= a534 + a533;
    a535 <= a535 + a534;
    a536 <= a536 + a535;
    a537 <= a537 + a536;
    a538 <= a538 + a537;
    a539 <= a539 + a538;
    a540 <= a540 + a539;
    a541 <= a541 + a540;
    a542 <= a542 + a541;
    a543 <= a543 + a542;
    a544 <= a544 + a543;
    a545 <= a545 + a544;
    a546 <= a546 + a545;
    a547 <= a547 + a546;
    a548 <= a548 + a547;
    a549 <= a549 + a548;
    a550 <= a550 + a549;
    a551 <= a551 + a550;
    a552 <= a552 + a551;
    a553 <= a553 + a552;
    a554 <= a554 + a553;
    a555 <= a555 + a554;
    a556 <= a556 + a555;
    a557 <= a557 + a556;
    a558 <= a558 + a557;
    a559 <= a559 + a558;
    a560 <= a560 + a559;
    a561 <= a561 + a560;
    a562 <= a562 + a561;
    a563 <= a563 + a562;
    a564 <= a564 + a563;
    a565 <= a565 + a564;
    a566 <= a566 + a565;
    a567 <= a567 + a566;
    a568 <= a568 + a567;
    a569 <= a569 + a568;
    a570 <= a570 + a569;
    a571 <= a571 + a570;
    a572 <= a572 + a571;
    a573 <= a573 + a572;
    a574 <= a574 + a573;
    a575 <= a575 + a574;
    a576 <= a576 + a575;
    a577 <= a577 + a576;
    a578 <= a578 + a577;
    a579 <= a579 + a578;
    a580 <= a580 + a579;
    a581 <= a581 + a580;
    a582 <= a582 + a581;
    a583 <= a583 + a582;
    a584 <= a584 + a583;
    a585 <= a585 + a584;
    a586 <= a586 + a585;
    a587 <= a587 + a586;
    a588 <= a588 + a587;
    a589 <= a589 + a588;
    a590 <= a590 + a589;
    a591 <= a591 + a590;
    a592 <= a592 + a591;
    a593 <= a593 + a592;
    a594 <= a594 + a593;
    a595 <= a595 + a594;
    a596 <= a596 + a595;
    a597 <= a597 + a596;
    a598 <= a598 + a597;
    a599 <= a599 + a598;
    a600 <= a600 + a599;
    a601 <= a601 + a600;
    a602 <= a602 + a601;
    a603 <= a603 + a602;
    a604 <= a604 + a603;
    a605 <= a605 + a604;
    a606 <= a606 + a605;
    a607 <= a607 + a606;
    a608 <= a608 + a607;
    a609 <= a609 + a608;
    a610 <= a610 + a609;
    a611 <= a611 + a610;
    a612 <= a612 + a611;
    a613 <= a613 + a612;
    a614 <= a614 + a613;
    a615 <= a615 + a614;
    a616 <= a616 + a615;
    a617 <= a617 + a616;
    a618 <= a618 + a617;
    a619 <= a619 + a618;
    a620 <= a620 + a619;
    a621 <= a621 + a620;
    a622 <= a622 + a621;
    a623 <= a623 + a622;
    a624 <= a624 + a623;
    a625 <= a625 + a624;
    a626 <= a626 + a625;
    a627 <= a627 + a626;
    a628 <= a628 + a627;
    a629 <= a629 + a628;
    a630 <= a630 + a629;
    a631 <= a631 + a630;
    a632 <= a632 + a631;
    a633 <= a633 + a632;
    a634 <= a634 + a633;
    a635 <= a635 + a634;
    a636 <= a636 + a635;
    a637 <= a637 + a636;
    a638 <= a638 + a637;
    a639 <= a639 + a638;
    a640 <= a640 + a639;
    a641 <= a641 + a640;
    a642 <= a642 + a641;
    a643 <= a643 + a642;
    a644 <= a644 + a643;
    a645 <= a645 + a644;
    a646 <= a646 + a645;
    a647 <= a647 + a646;
    a648 <= a648 + a647;
    a649 <= a649 + a648;
    a650 <= a650 + a649;
    a651 <= a651 + a650;
    a652 <= a652 + a651;
    a653 <= a653 + a652;
    a654 <= a654 + a653;
    a655 <= a655 + a654;
    a656 <= a656 + a655;
    a657 <= a657 + a656;
    a658 <= a658 + a657;
    a659 <= a659 + a658;
    a660 <= a660 + a659;
    a661 <= a661 + a660;
    a662 <= a662 + a661;
    a663 <= a663 + a662;
    a664 <= a664 + a663;
    a665 <= a665 + a664;
    a666 <= a666 + a665;
    a667 <= a667 + a666;
    a668 <= a668 + a667;
    a669 <= a669 + a668;
    a670 <= a670 + a669;
    a671 <= a671 + a670;
    a672 <= a672 + a671;
    a673 <= a673 + a672;
    a674 <= a674 + a673;
    a675 <= a675 + a674;
    a676 <= a676 + a675;
    a677 <= a677 + a676;
    a678 <= a678 + a677;
    a679 <= a679 + a678;
    a680 <= a680 + a679;
    a681 <= a681 + a680;
    a682 <= a682 + a681;
    a683 <= a683 + a682;
    a684 <= a684 + a683;
    a685 <= a685 + a684;
    a686 <= a686 + a685;
    a687 <= a687 + a686;
    a688 <= a688 + a687;
    a689 <= a689 + a688;
    a690 <= a690 + a689;
    a691 <= a691 + a690;
    a692 <= a692 + a691;
    a693 <= a693 + a692;
    a694 <= a694 + a693;
    a695 <= a695 + a694;
    a696 <= a696 + a695;
    a697 <= a697 + a696;
    a698 <= a698 + a697;
    a699 <= a699 + a698;
    a700 <= a700 + a699;
    a701 <= a701 + a700;
    a702 <= a702 + a701;
    a703 <= a703 + a702;
    a704 <= a704 + a703;
    a705 <= a705 + a704;
    a706 <= a706 + a705;
    a707 <= a707 + a706;
    a708 <= a708 + a707;
    a709 <= a709 + a708;
    a710 <= a710 + a709;
    a711 <= a711 + a710;
    a712 <= a712 + a711;
    a713 <= a713 + a712;
    a714 <= a714 + a713;
    a715 <= a715 + a714;
    a716 <= a716 + a715;
    a717 <= a717 + a716;
    a718 <= a718 + a717;
    a719 <= a719 + a718;
    a720 <= a720 + a719;
    a721 <= a721 + a720;
    a722 <= a722 + a721;
    a723 <= a723 + a722;
    a724 <= a724 + a723;
    a725 <= a725 + a724;
    a726 <= a726 + a725;
    a727 <= a727 + a726;
    a728 <= a728 + a727;
    a729 <= a729 + a728;
    a730 <= a730 + a729;
    a731 <= a731 + a730;
    a732 <= a732 + a731;
    a733 <= a733 + a732;
    a734 <= a734 + a733;
    a735 <= a735 + a734;
    a736 <= a736 + a735;
    a737 <= a737 + a736;
    a738 <= a738 + a737;
    a739 <= a739 + a738;
    a740 <= a740 + a739;
    a741 <= a741 + a740;
    a742 <= a742 + a741;
    a743 <= a743 + a742;
    a744 <= a744 + a743;
    a745 <= a745 + a744;
    a746 <= a746 + a745;
    a747 <= a747 + a746;
    a748 <= a748 + a747;
    a749 <= a749 + a748;
    a750 <= a750 + a749;
    a751 <= a751 + a750;
    a752 <= a752 + a751;
    a753 <= a753 + a752;
    a754 <= a754 + a753;
    a755 <= a755 + a754;
    a756 <= a756 + a755;
    a757 <= a757 + a756;
    a758 <= a758 + a757;
    a759 <= a759 + a758;
    a760 <= a760 + a759;
    a761 <= a761 + a760;
    a762 <= a762 + a761;
    a763 <= a763 + a762;
    a764 <= a764 + a763;
    a765 <= a765 + a764;
    a766 <= a766 + a765;
    a767 <= a767 + a766;
    a768 <= a768 + a767;
    a769 <= a769 + a768;
    a770 <= a770 + a769;
    a771 <= a771 + a770;
    a772 <= a772 + a771;
    a773 <= a773 + a772;
    a774 <= a774 + a773;
    a775 <= a775 + a774;
    a776 <= a776 + a775;
    a777 <= a777 + a776;
    a778 <= a778 + a777;
    a779 <= a779 + a778;
    a780 <= a780 + a779;
    a781 <= a781 + a780;
    a782 <= a782 + a781;
    a783 <= a783 + a782;
    a784 <= a784 + a783;
    a785 <= a785 + a784;
    a786 <= a786 + a785;
    a787 <= a787 + a786;
    a788 <= a788 + a787;
    a789 <= a789 + a788;
    a790 <= a790 + a789;
    a791 <= a791 + a790;
    a792 <= a792 + a791;
    a793 <= a793 + a792;
    a794 <= a794 + a793;
    a795 <= a795 + a794;
    a796 <= a796 + a795;
    a797 <= a797 + a796;
    a798 <= a798 + a797;
    a799 <= a799 + a798;
    a800 <= a800 + a799;
    a801 <= a801 + a800;
    a802 <= a802 + a801;
    a803 <= a803 + a802;
    a804 <= a804 + a803;
    a805 <= a805 + a804;
    a806 <= a806 + a805;
    a807 <= a807 + a806;
    a808 <= a808 + a807;
    a809 <= a809 + a808;
    a810 <= a810 + a809;
    a811 <= a811 + a810;
    a812 <= a812 + a811;
    a813 <= a813 + a812;
    a814 <= a814 + a813;
    a815 <= a815 + a814;
    a816 <= a816 + a815;
    a817 <= a817 + a816;
    a818 <= a818 + a817;
    a819 <= a819 + a818;
    a820 <= a820 + a819;
    a821 <= a821 + a820;
    a822 <= a822 + a821;
    a823 <= a823 + a822;
    a824 <= a824 + a823;
    a825 <= a825 + a824;
    a826 <= a826 + a825;
    a827 <= a827 + a826;
    a828 <= a828 + a827;
    a829 <= a829 + a828;
    a830 <= a830 + a829;
    a831 <= a831 + a830;
    a832 <= a832 + a831;
    a833 <= a833 + a832;
    a834 <= a834 + a833;
    a835 <= a835 + a834;
    a836 <= a836 + a835;
    a837 <= a837 + a836;
    a838 <= a838 + a837;
    a839 <= a839 + a838;
    a840 <= a840 + a839;
    a841 <= a841 + a840;
    a842 <= a842 + a841;
    a843 <= a843 + a842;
    a844 <= a844 + a843;
    a845 <= a845 + a844;
    a846 <= a846 + a845;
    a847 <= a847 + a846;
    a848 <= a848 + a847;
    a849 <= a849 + a848;
    a850 <= a850 + a849;
    a851 <= a851 + a850;
    a852 <= a852 + a851;
    a853 <= a853 + a852;
    a854 <= a854 + a853;
    a855 <= a855 + a854;
    a856 <= a856 + a855;
    a857 <= a857 + a856;
    a858 <= a858 + a857;
    a859 <= a859 + a858;
    a860 <= a860 + a859;
    a861 <= a861 + a860;
    a862 <= a862 + a861;
    a863 <= a863 + a862;
    a864 <= a864 + a863;
    a865 <= a865 + a864;
    a866 <= a866 + a865;
    a867 <= a867 + a866;
    a868 <= a868 + a867;
    a869 <= a869 + a868;
    a870 <= a870 + a869;
    a871 <= a871 + a870;
    a872 <= a872 + a871;
    a873 <= a873 + a872;
    a874 <= a874 + a873;
    a875 <= a875 + a874;
    a876 <= a876 + a875;
    a877 <= a877 + a876;
    a878 <= a878 + a877;
    a879 <= a879 + a878;
    a880 <= a880 + a879;
    a881 <= a881 + a880;
    a882 <= a882 + a881;
    a883 <= a883 + a882;
    a884 <= a884 + a883;
    a885 <= a885 + a884;
    a886 <= a886 + a885;
    a887 <= a887 + a886;
    a888 <= a888 + a887;
    a889 <= a889 + a888;
    a890 <= a890 + a889;
    a891 <= a891 + a890;
    a892 <= a892 + a891;
    a893 <= a893 + a892;
    a894 <= a894 + a893;
    a895 <= a895 + a894;
    a896 <= a896 + a895;
    a897 <= a897 + a896;
    a898 <= a898 + a897;
    a899 <= a899 + a898;
    a900 <= a900 + a899;
    a901 <= a901 + a900;
    a902 <= a902 + a901;
    a903 <= a903 + a902;
    a904 <= a904 + a903;
    a905 <= a905 + a904;
    a906 <= a906 + a905;
    a907 <= a907 + a906;
    a908 <= a908 + a907;
    a909 <= a909 + a908;
    a910 <= a910 + a909;
    a911 <= a911 + a910;
    a912 <= a912 + a911;
    a913 <= a913 + a912;
    a914 <= a914 + a913;
    a915 <= a915 + a914;
    a916 <= a916 + a915;
    a917 <= a917 + a916;
    a918 <= a918 + a917;
    a919 <= a919 + a918;
    a920 <= a920 + a919;
    a921 <= a921 + a920;
    a922 <= a922 + a921;
    a923 <= a923 + a922;
    a924 <= a924 + a923;
    a925 <= a925 + a924;
    a926 <= a926 + a925;
    a927 <= a927 + a926;
    a928 <= a928 + a927;
    a929 <= a929 + a928;
    a930 <= a930 + a929;
    a931 <= a931 + a930;
    a932 <= a932 + a931;
    a933 <= a933 + a932;
    a934 <= a934 + a933;
    a935 <= a935 + a934;
    a936 <= a936 + a935;
    a937 <= a937 + a936;
    a938 <= a938 + a937;
    a939 <= a939 + a938;
    a940 <= a940 + a939;
    a941 <= a941 + a940;
    a942 <= a942 + a941;
    a943 <= a943 + a942;
    a944 <= a944 + a943;
    a945 <= a945 + a944;
    a946 <= a946 + a945;
    a947 <= a947 + a946;
    a948 <= a948 + a947;
    a949 <= a949 + a948;
    a950 <= a950 + a949;
    a951 <= a951 + a950;
    a952 <= a952 + a951;
    a953 <= a953 + a952;
    a954 <= a954 + a953;
    a955 <= a955 + a954;
    a956 <= a956 + a955;
    a957 <= a957 + a956;
    a958 <= a958 + a957;
    a959 <= a959 + a958;
    a960 <= a960 + a959;
    a961 <= a961 + a960;
    a962 <= a962 + a961;
    a963 <= a963 + a962;
    a964 <= a964 + a963;
    a965 <= a965 + a964;
    a966 <= a966 + a965;
    a967 <= a967 + a966;
    a968 <= a968 + a967;
    a969 <= a969 + a968;
    a970 <= a970 + a969;
    a971 <= a971 + a970;
    a972 <= a972 + a971;
    a973 <= a973 + a972;
    a974 <= a974 + a973;
    a975 <= a975 + a974;
    a976 <= a976 + a975;
    a977 <= a977 + a976;
    a978 <= a978 + a977;
    a979 <= a979 + a978;
    a980 <= a980 + a979;
    a981 <= a981 + a980;
    a982 <= a982 + a981;
    a983 <= a983 + a982;
    a984 <= a984 + a983;
    a985 <= a985 + a984;
    a986 <= a986 + a985;
    a987 <= a987 + a986;
    a988 <= a988 + a987;
    a989 <= a989 + a988;
    a990 <= a990 + a989;
    a991 <= a991 + a990;
    a992 <= a992 + a991;
    a993 <= a993 + a992;
    a994 <= a994 + a993;
    a995 <= a995 + a994;
    a996 <= a996 + a995;
    a997 <= a997 + a996;
    a998 <= a998 + a997;
    a999 <= a999 + a998;
    a1000 <= a1000 + a999;
    a1001 <= a1001 + a1000;
    a1002 <= a1002 + a1001;
    a1003 <= a1003 + a1002;
    a1004 <= a1004 + a1003;
    a1005 <= a1005 + a1004;
    a1006 <= a1006 + a1005;
    a1007 <= a1007 + a1006;
    a1008 <= a1008 + a1007;
    a1009 <= a1009 + a1008;
    a1010 <= a1010 + a1009;
    a1011 <= a1011 + a1010;
    a1012 <= a1012 + a1011;
    a1013 <= a1013 + a1012;
    a1014 <= a1014 + a1013;
    a1015 <= a1015 + a1014;
    a1016 <= a1016 + a1015;
    a1017 <= a1017 + a1016;
    a1018 <= a1018 + a1017;
    a1019 <= a1019 + a1018;
    a1020 <= a1020 + a1019;
    a1021 <= a1021 + a1020;
    a1022 <= a1022 + a1021;
    a1023 <= a1023 + a1022;
    a1024 <= a1024 + a1023;
    a1025 <= a1025 + a1024;
    a1026 <= a1026 + a1025;
    a1027 <= a1027 + a1026;
    a1028 <= a1028 + a1027;
    a1029 <= a1029 + a1028;
    a1030 <= a1030 + a1029;
    a1031 <= a1031 + a1030;
    a1032 <= a1032 + a1031;
    a1033 <= a1033 + a1032;
    a1034 <= a1034 + a1033;
    a1035 <= a1035 + a1034;
    a1036 <= a1036 + a1035;
    a1037 <= a1037 + a1036;
    a1038 <= a1038 + a1037;
    a1039 <= a1039 + a1038;
    a1040 <= a1040 + a1039;
    a1041 <= a1041 + a1040;
    a1042 <= a1042 + a1041;
    a1043 <= a1043 + a1042;
    a1044 <= a1044 + a1043;
    a1045 <= a1045 + a1044;
    a1046 <= a1046 + a1045;
    a1047 <= a1047 + a1046;
    a1048 <= a1048 + a1047;
    a1049 <= a1049 + a1048;
    a1050 <= a1050 + a1049;
    a1051 <= a1051 + a1050;
    a1052 <= a1052 + a1051;
    a1053 <= a1053 + a1052;
    a1054 <= a1054 + a1053;
    a1055 <= a1055 + a1054;
    a1056 <= a1056 + a1055;
    a1057 <= a1057 + a1056;
    a1058 <= a1058 + a1057;
    a1059 <= a1059 + a1058;
    a1060 <= a1060 + a1059;
    a1061 <= a1061 + a1060;
    a1062 <= a1062 + a1061;
    a1063 <= a1063 + a1062;
    a1064 <= a1064 + a1063;
    a1065 <= a1065 + a1064;
    a1066 <= a1066 + a1065;
    a1067 <= a1067 + a1066;
    a1068 <= a1068 + a1067;
    a1069 <= a1069 + a1068;
    a1070 <= a1070 + a1069;
    a1071 <= a1071 + a1070;
    a1072 <= a1072 + a1071;
    a1073 <= a1073 + a1072;
    a1074 <= a1074 + a1073;
    a1075 <= a1075 + a1074;
    a1076 <= a1076 + a1075;
    a1077 <= a1077 + a1076;
    a1078 <= a1078 + a1077;
    a1079 <= a1079 + a1078;
    a1080 <= a1080 + a1079;
    a1081 <= a1081 + a1080;
    a1082 <= a1082 + a1081;
    a1083 <= a1083 + a1082;
    a1084 <= a1084 + a1083;
    a1085 <= a1085 + a1084;
    a1086 <= a1086 + a1085;
    a1087 <= a1087 + a1086;
    a1088 <= a1088 + a1087;
    a1089 <= a1089 + a1088;
    a1090 <= a1090 + a1089;
    a1091 <= a1091 + a1090;
    a1092 <= a1092 + a1091;
    a1093 <= a1093 + a1092;
    a1094 <= a1094 + a1093;
    a1095 <= a1095 + a1094;
    a1096 <= a1096 + a1095;
    a1097 <= a1097 + a1096;
    a1098 <= a1098 + a1097;
    a1099 <= a1099 + a1098;
    a1100 <= a1100 + a1099;
    a1101 <= a1101 + a1100;
    a1102 <= a1102 + a1101;
    a1103 <= a1103 + a1102;
    a1104 <= a1104 + a1103;
    a1105 <= a1105 + a1104;
    a1106 <= a1106 + a1105;
    a1107 <= a1107 + a1106;
    a1108 <= a1108 + a1107;
    a1109 <= a1109 + a1108;
    a1110 <= a1110 + a1109;
    a1111 <= a1111 + a1110;
    a1112 <= a1112 + a1111;
    a1113 <= a1113 + a1112;
    a1114 <= a1114 + a1113;
    a1115 <= a1115 + a1114;
    a1116 <= a1116 + a1115;
    a1117 <= a1117 + a1116;
    a1118 <= a1118 + a1117;
    a1119 <= a1119 + a1118;
    a1120 <= a1120 + a1119;
    a1121 <= a1121 + a1120;
    a1122 <= a1122 + a1121;
    a1123 <= a1123 + a1122;
    a1124 <= a1124 + a1123;
    a1125 <= a1125 + a1124;
    a1126 <= a1126 + a1125;
    a1127 <= a1127 + a1126;
    a1128 <= a1128 + a1127;
    a1129 <= a1129 + a1128;
    a1130 <= a1130 + a1129;
    a1131 <= a1131 + a1130;
    a1132 <= a1132 + a1131;
    a1133 <= a1133 + a1132;
    a1134 <= a1134 + a1133;
    a1135 <= a1135 + a1134;
    a1136 <= a1136 + a1135;
    a1137 <= a1137 + a1136;
    a1138 <= a1138 + a1137;
    a1139 <= a1139 + a1138;
    a1140 <= a1140 + a1139;
    a1141 <= a1141 + a1140;
    a1142 <= a1142 + a1141;
    a1143 <= a1143 + a1142;
    a1144 <= a1144 + a1143;
    a1145 <= a1145 + a1144;
    a1146 <= a1146 + a1145;
    a1147 <= a1147 + a1146;
    a1148 <= a1148 + a1147;
    a1149 <= a1149 + a1148;
    a1150 <= a1150 + a1149;
    a1151 <= a1151 + a1150;
    a1152 <= a1152 + a1151;
    a1153 <= a1153 + a1152;
    a1154 <= a1154 + a1153;
    a1155 <= a1155 + a1154;
    a1156 <= a1156 + a1155;
    a1157 <= a1157 + a1156;
    a1158 <= a1158 + a1157;
    a1159 <= a1159 + a1158;
    a1160 <= a1160 + a1159;
    a1161 <= a1161 + a1160;
    a1162 <= a1162 + a1161;
    a1163 <= a1163 + a1162;
    a1164 <= a1164 + a1163;
    a1165 <= a1165 + a1164;
    a1166 <= a1166 + a1165;
    a1167 <= a1167 + a1166;
    a1168 <= a1168 + a1167;
    a1169 <= a1169 + a1168;
    a1170 <= a1170 + a1169;
    a1171 <= a1171 + a1170;
    a1172 <= a1172 + a1171;
    a1173 <= a1173 + a1172;
    a1174 <= a1174 + a1173;
    a1175 <= a1175 + a1174;
    a1176 <= a1176 + a1175;
    a1177 <= a1177 + a1176;
    a1178 <= a1178 + a1177;
    a1179 <= a1179 + a1178;
    a1180 <= a1180 + a1179;
    a1181 <= a1181 + a1180;
    a1182 <= a1182 + a1181;
    a1183 <= a1183 + a1182;
    a1184 <= a1184 + a1183;
    a1185 <= a1185 + a1184;
    a1186 <= a1186 + a1185;
    a1187 <= a1187 + a1186;
    a1188 <= a1188 + a1187;
    a1189 <= a1189 + a1188;
    a1190 <= a1190 + a1189;
    a1191 <= a1191 + a1190;
    a1192 <= a1192 + a1191;
    a1193 <= a1193 + a1192;
    a1194 <= a1194 + a1193;
    a1195 <= a1195 + a1194;
    a1196 <= a1196 + a1195;
    a1197 <= a1197 + a1196;
    a1198 <= a1198 + a1197;
    a1199 <= a1199 + a1198;
    a1200 <= a1200 + a1199;
    a1201 <= a1201 + a1200;
    a1202 <= a1202 + a1201;
    a1203 <= a1203 + a1202;
    a1204 <= a1204 + a1203;
    a1205 <= a1205 + a1204;
    a1206 <= a1206 + a1205;
    a1207 <= a1207 + a1206;
    a1208 <= a1208 + a1207;
    a1209 <= a1209 + a1208;
    a1210 <= a1210 + a1209;
    a1211 <= a1211 + a1210;
    a1212 <= a1212 + a1211;
    a1213 <= a1213 + a1212;
    a1214 <= a1214 + a1213;
    a1215 <= a1215 + a1214;
    a1216 <= a1216 + a1215;
    a1217 <= a1217 + a1216;
    a1218 <= a1218 + a1217;
    a1219 <= a1219 + a1218;
    a1220 <= a1220 + a1219;
    a1221 <= a1221 + a1220;
    a1222 <= a1222 + a1221;
    a1223 <= a1223 + a1222;
    a1224 <= a1224 + a1223;
    a1225 <= a1225 + a1224;
    a1226 <= a1226 + a1225;
    a1227 <= a1227 + a1226;
    a1228 <= a1228 + a1227;
    a1229 <= a1229 + a1228;
    a1230 <= a1230 + a1229;
    a1231 <= a1231 + a1230;
    a1232 <= a1232 + a1231;
    a1233 <= a1233 + a1232;
    a1234 <= a1234 + a1233;
    a1235 <= a1235 + a1234;
    a1236 <= a1236 + a1235;
    a1237 <= a1237 + a1236;
    a1238 <= a1238 + a1237;
    a1239 <= a1239 + a1238;
    a1240 <= a1240 + a1239;
    a1241 <= a1241 + a1240;
    a1242 <= a1242 + a1241;
    a1243 <= a1243 + a1242;
    a1244 <= a1244 + a1243;
    a1245 <= a1245 + a1244;
    a1246 <= a1246 + a1245;
    a1247 <= a1247 + a1246;
    a1248 <= a1248 + a1247;
    a1249 <= a1249 + a1248;
    a1250 <= a1250 + a1249;
    a1251 <= a1251 + a1250;
    a1252 <= a1252 + a1251;
    a1253 <= a1253 + a1252;
    a1254 <= a1254 + a1253;
    a1255 <= a1255 + a1254;
    a1256 <= a1256 + a1255;
    a1257 <= a1257 + a1256;
    a1258 <= a1258 + a1257;
    a1259 <= a1259 + a1258;
    a1260 <= a1260 + a1259;
    a1261 <= a1261 + a1260;
    a1262 <= a1262 + a1261;
    a1263 <= a1263 + a1262;
    a1264 <= a1264 + a1263;
    a1265 <= a1265 + a1264;
    a1266 <= a1266 + a1265;
    a1267 <= a1267 + a1266;
    a1268 <= a1268 + a1267;
    a1269 <= a1269 + a1268;
    a1270 <= a1270 + a1269;
    a1271 <= a1271 + a1270;
    a1272 <= a1272 + a1271;
    a1273 <= a1273 + a1272;
    a1274 <= a1274 + a1273;
    a1275 <= a1275 + a1274;
    a1276 <= a1276 + a1275;
    a1277 <= a1277 + a1276;
    a1278 <= a1278 + a1277;
    a1279 <= a1279 + a1278;
    a1280 <= a1280 + a1279;
    a1281 <= a1281 + a1280;
    a1282 <= a1282 + a1281;
    a1283 <= a1283 + a1282;
    a1284 <= a1284 + a1283;
    a1285 <= a1285 + a1284;
    a1286 <= a1286 + a1285;
    a1287 <= a1287 + a1286;
    a1288 <= a1288 + a1287;
    a1289 <= a1289 + a1288;
    a1290 <= a1290 + a1289;
    a1291 <= a1291 + a1290;
    a1292 <= a1292 + a1291;
    a1293 <= a1293 + a1292;
    a1294 <= a1294 + a1293;
    a1295 <= a1295 + a1294;
    a1296 <= a1296 + a1295;
    a1297 <= a1297 + a1296;
    a1298 <= a1298 + a1297;
    a1299 <= a1299 + a1298;
    a1300 <= a1300 + a1299;
    a1301 <= a1301 + a1300;
    a1302 <= a1302 + a1301;
    a1303 <= a1303 + a1302;
    a1304 <= a1304 + a1303;
    a1305 <= a1305 + a1304;
    a1306 <= a1306 + a1305;
    a1307 <= a1307 + a1306;
    a1308 <= a1308 + a1307;
    a1309 <= a1309 + a1308;
    a1310 <= a1310 + a1309;
    a1311 <= a1311 + a1310;
    a1312 <= a1312 + a1311;
    a1313 <= a1313 + a1312;
    a1314 <= a1314 + a1313;
    a1315 <= a1315 + a1314;
    a1316 <= a1316 + a1315;
    a1317 <= a1317 + a1316;
    a1318 <= a1318 + a1317;
    a1319 <= a1319 + a1318;
    a1320 <= a1320 + a1319;
    a1321 <= a1321 + a1320;
    a1322 <= a1322 + a1321;
    a1323 <= a1323 + a1322;
    a1324 <= a1324 + a1323;
    a1325 <= a1325 + a1324;
    a1326 <= a1326 + a1325;
    a1327 <= a1327 + a1326;
    a1328 <= a1328 + a1327;
    a1329 <= a1329 + a1328;
    a1330 <= a1330 + a1329;
    a1331 <= a1331 + a1330;
    a1332 <= a1332 + a1331;
    a1333 <= a1333 + a1332;
    a1334 <= a1334 + a1333;
    a1335 <= a1335 + a1334;
    a1336 <= a1336 + a1335;
    a1337 <= a1337 + a1336;
    a1338 <= a1338 + a1337;
    a1339 <= a1339 + a1338;
    a1340 <= a1340 + a1339;
    a1341 <= a1341 + a1340;
    a1342 <= a1342 + a1341;
    a1343 <= a1343 + a1342;
    a1344 <= a1344 + a1343;
    a1345 <= a1345 + a1344;
    a1346 <= a1346 + a1345;
    a1347 <= a1347 + a1346;
    a1348 <= a1348 + a1347;
    a1349 <= a1349 + a1348;
    a1350 <= a1350 + a1349;
    a1351 <= a1351 + a1350;
    a1352 <= a1352 + a1351;
    a1353 <= a1353 + a1352;
    a1354 <= a1354 + a1353;
    a1355 <= a1355 + a1354;
    a1356 <= a1356 + a1355;
    a1357 <= a1357 + a1356;
    a1358 <= a1358 + a1357;
    a1359 <= a1359 + a1358;
    a1360 <= a1360 + a1359;
    a1361 <= a1361 + a1360;
    a1362 <= a1362 + a1361;
    a1363 <= a1363 + a1362;
    a1364 <= a1364 + a1363;
    a1365 <= a1365 + a1364;
    a1366 <= a1366 + a1365;
    a1367 <= a1367 + a1366;
    a1368 <= a1368 + a1367;
    a1369 <= a1369 + a1368;
    a1370 <= a1370 + a1369;
    a1371 <= a1371 + a1370;
    a1372 <= a1372 + a1371;
    a1373 <= a1373 + a1372;
    a1374 <= a1374 + a1373;
    a1375 <= a1375 + a1374;
    a1376 <= a1376 + a1375;
    a1377 <= a1377 + a1376;
    a1378 <= a1378 + a1377;
    a1379 <= a1379 + a1378;
    a1380 <= a1380 + a1379;
    a1381 <= a1381 + a1380;
    a1382 <= a1382 + a1381;
    a1383 <= a1383 + a1382;
    a1384 <= a1384 + a1383;
    a1385 <= a1385 + a1384;
    a1386 <= a1386 + a1385;
    a1387 <= a1387 + a1386;
    a1388 <= a1388 + a1387;
    a1389 <= a1389 + a1388;
    a1390 <= a1390 + a1389;
    a1391 <= a1391 + a1390;
    a1392 <= a1392 + a1391;
    a1393 <= a1393 + a1392;
    a1394 <= a1394 + a1393;
    a1395 <= a1395 + a1394;
    a1396 <= a1396 + a1395;
    a1397 <= a1397 + a1396;
    a1398 <= a1398 + a1397;
    a1399 <= a1399 + a1398;
    a1400 <= a1400 + a1399;
    a1401 <= a1401 + a1400;
    a1402 <= a1402 + a1401;
    a1403 <= a1403 + a1402;
    a1404 <= a1404 + a1403;
    a1405 <= a1405 + a1404;
    a1406 <= a1406 + a1405;
    a1407 <= a1407 + a1406;
    a1408 <= a1408 + a1407;
    a1409 <= a1409 + a1408;
    a1410 <= a1410 + a1409;
    a1411 <= a1411 + a1410;
    a1412 <= a1412 + a1411;
    a1413 <= a1413 + a1412;
    a1414 <= a1414 + a1413;
    a1415 <= a1415 + a1414;
    a1416 <= a1416 + a1415;
    a1417 <= a1417 + a1416;
    a1418 <= a1418 + a1417;
    a1419 <= a1419 + a1418;
    a1420 <= a1420 + a1419;
    a1421 <= a1421 + a1420;
    a1422 <= a1422 + a1421;
    a1423 <= a1423 + a1422;
    a1424 <= a1424 + a1423;
    a1425 <= a1425 + a1424;
    a1426 <= a1426 + a1425;
    a1427 <= a1427 + a1426;
    a1428 <= a1428 + a1427;
    a1429 <= a1429 + a1428;
    a1430 <= a1430 + a1429;
    a1431 <= a1431 + a1430;
    a1432 <= a1432 + a1431;
    a1433 <= a1433 + a1432;
    a1434 <= a1434 + a1433;
    a1435 <= a1435 + a1434;
    a1436 <= a1436 + a1435;
    a1437 <= a1437 + a1436;
    a1438 <= a1438 + a1437;
    a1439 <= a1439 + a1438;
    a1440 <= a1440 + a1439;
    a1441 <= a1441 + a1440;
    a1442 <= a1442 + a1441;
    a1443 <= a1443 + a1442;
    a1444 <= a1444 + a1443;
    a1445 <= a1445 + a1444;
    a1446 <= a1446 + a1445;
    a1447 <= a1447 + a1446;
    a1448 <= a1448 + a1447;
    a1449 <= a1449 + a1448;
    a1450 <= a1450 + a1449;
    a1451 <= a1451 + a1450;
    a1452 <= a1452 + a1451;
    a1453 <= a1453 + a1452;
    a1454 <= a1454 + a1453;
    a1455 <= a1455 + a1454;
    a1456 <= a1456 + a1455;
    a1457 <= a1457 + a1456;
    a1458 <= a1458 + a1457;
    a1459 <= a1459 + a1458;
    a1460 <= a1460 + a1459;
    a1461 <= a1461 + a1460;
    a1462 <= a1462 + a1461;
    a1463 <= a1463 + a1462;
    a1464 <= a1464 + a1463;
    a1465 <= a1465 + a1464;
    a1466 <= a1466 + a1465;
    a1467 <= a1467 + a1466;
    a1468 <= a1468 + a1467;
    a1469 <= a1469 + a1468;
    a1470 <= a1470 + a1469;
    a1471 <= a1471 + a1470;
    a1472 <= a1472 + a1471;
    a1473 <= a1473 + a1472;
    a1474 <= a1474 + a1473;
    a1475 <= a1475 + a1474;
    a1476 <= a1476 + a1475;
    a1477 <= a1477 + a1476;
    a1478 <= a1478 + a1477;
    a1479 <= a1479 + a1478;
    a1480 <= a1480 + a1479;
    a1481 <= a1481 + a1480;
    a1482 <= a1482 + a1481;
    a1483 <= a1483 + a1482;
    a1484 <= a1484 + a1483;
    a1485 <= a1485 + a1484;
    a1486 <= a1486 + a1485;
    a1487 <= a1487 + a1486;
    a1488 <= a1488 + a1487;
    a1489 <= a1489 + a1488;
    a1490 <= a1490 + a1489;
    a1491 <= a1491 + a1490;
    a1492 <= a1492 + a1491;
    a1493 <= a1493 + a1492;
    a1494 <= a1494 + a1493;
    a1495 <= a1495 + a1494;
    a1496 <= a1496 + a1495;
    a1497 <= a1497 + a1496;
    a1498 <= a1498 + a1497;
    a1499 <= a1499 + a1498;
    a1500 <= a1500 + a1499;
  end

endmodule
